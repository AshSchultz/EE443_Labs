-- LIBRARY ieee;
-- USE ieee.std_logic_1164.all;

-- entity sim_REG8 is
-- end entity sim_REG8;
-- architecture Behavioral of sim_REG8 is
    
--     SIGNAL X, Y : std_logic_vector := '0';
--     SIGNAL E, C : std_logic := '0';

-- begin
    
--     dut : entity work.half_adder
--         port map(
--             x => X,
--             EN =>
--             CLK : in std_logic;
--             y : out std_logic_vector(7 downto 0)
--         );
--     end entity REG8;
    
-- end architecture Behavioral;